library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity datapath is

end entity;

architecture basic of datapath is

begin
end basic;