library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IRMux is 

port(
		instr: in std_logic_vector(15 downto 0);
		
	);

end entity;

architecture basic of IRMux is

begin

end basic;